module muxdisplay(
input [7:0] E0,
input [7:0] E1,
input Escolha,
output [7:0]Saida
);


endmodule